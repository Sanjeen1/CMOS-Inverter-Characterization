.include ./tsmc180.txt

m0 out in Gnd 0 nfet l=0.2u w =10u
m1 out in Vdd vdd pfet l=0.4u w= 10u
cl out Gnd 1p

Vdd vdd Gnd 1.8
Vdin in Gnd pulse(0 1.8 1p 10p 10p 10n 20n)

.control
foreach width 1u 10u 20u 100u

alter m1 w = $width

dc vdin 0 1.8 0.1m

meas dc Vm find v(in) when v(out)=v(in)
print Vm    
end
.endc
.end