.include ./tsmc180.txt

m0 out in Gnd 0 nfet l=0.2u w = 10u
m1 out in Vdd vdd pfet l=0.4u w= 10u
cl out Gnd 1f

Vdd vdd Gnd 1.8
Vdin in Gnd pulse(0 1.8 1p 10p 10p 10n 20n)

.dc Vdin 0 1.8 0.01
.control
foreach width 10u 20u 30u

alter m1 w = $width
 
run

set color0=white
set color1=black
set color2=red
set color3=blue
set color4=green
set xbrushwidth=3
end
plot dc1.out dc2.out dc3.out vs in title 'Pmos width vary'

.endc
.end


