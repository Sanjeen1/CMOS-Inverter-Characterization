.include ./tsmc180.txt

m0 out in Gnd 0 nfet l=0.2u w =10u
m1 out in Vdd vdd pfet l=0.4u w= 10u
cl out Gnd 1p

Vdd vdd Gnd 1.8
Vdin in Gnd pulse(0 1.8 1p 10p 10p 10n 20n)

.control
foreach width 1u 10u 20u

alter m1 w = $width

tran 10n 100n

let p = 1.8*(-Vdd#branch)
meas tran energy integ p from=0n to=20n
let power = energy/20n
print power

end
.endc
.end