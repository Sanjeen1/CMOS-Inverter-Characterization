* SPICE3 file created from (UNNAMED).ext - technology: tsmc

.include ./tsmc180.txt
.option scale=0.06u


Vdd vdd Gnd 1.8
Vdin in Gnd pulse(0 1.8 1p 10p 10p 10n 20n)





M1000 out in Gnd Gnd nfet w=9 l=3
+  ad=143 pd=50 as=90 ps=38
M1001 out in vdd vdd pfet w=8 l=3
+  ad=128 pd=48 as=80 ps=36

.control
run
setplot tran
plot out  in+8


set color0=white
set color1=black
set color2=red
set color3=blue
set xbrushwidth=3


.endc

.tran 10n 100n 
.measure tran T_rise trig v(out) val = 0.1*vdd rise = 1 targ v(out) val = 0.9*vdd rise = 1
.measure tran T_fall trig v(out) val = 0.9*vdd fall = 1 targ v(out) val = 0.1*vdd fall = 1
.measure tran T_delay trig v(in) val = 0.5*vdd rise = 1 targ v(out) val = 0.5*vdd rise = 1
.measure tran TPHL    trig v(in) val= 0.5*vdd  fall=1 targ v(out) val=0.5*vdd   rise=1
.measure tran TPLH   trig v(in) val=0.5*vdd   rise=1 targ v(out) val=0.5*vdd fall=1

                 
                 

                 
.end

