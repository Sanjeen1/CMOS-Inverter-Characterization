.include ./tsmc180.txt

m0 out in Gnd 0 nfet l=0.2u w =10u
m1 out in Vdd vdd pfet l=0.4u w= 10u
cl out Gnd 1p

Vdd vdd Gnd 1.8
Vdin in Gnd pulse(0 1.8 1p 10p 10p 10n 20n)

.control
foreach width 1u 10u 20u

alter m1 w = $width

tran 10n 100n

meas tran vd_max MAX v(out) from=0.1n to =5n
meas tran vd_min MIN v(out) from=1n to =10n

let low = vd_min + 0.1*(vd_max-vd_min)
let high = vd_min + 0.9*(vd_max - vd_min)

meas tran rise_t TRIG V(out) VAL=low rise=1 TARG V(out) VAL=high rise=1
meas tran fall_t TRIG V(out) VAL=high fall=1 TARG V(out) VAL=low fall=1

let mid = 0.5*(vd_min+vd_max)

meas tran tphl trig in val=0.9 rise=1 targ v(out) val=mid fall=1
meas tran tplh trig in val=0.9 fall=1 targ v(out) val=mid rise=1

let prop_delay = (tphl+tplh)/2
print prop_delay

end
.endc
.end